----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    03:28:46 03/25/2022 
-- Design Name: 
-- Module Name:    myDataTypes - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

package myDataTypes is
 
type array32 	is array (31 downto 0) 	of STD_LOGIC_VECTOR (31 downto 0);
   
end package ;
 


