
use IEEE.STD_LOGIC_1164.ALL;



entity FORWARN_UNIT is
end FORWARN_UNIT;

architecture Behavioral of FORWARN_UNIT is

begin


end Behavioral;

